library ieee;
use ieee.std_logic_1164.all;

entity uROM is
port(
	ADD: in std_logic_vector(3 downto 0);
	Q: out std_logic_vector(45 downto 0)
);
end entity;

architecture behavioral of uROM is

begin
process(ADD)
begin
	case ADD is
     	when "0000" => Q <= "0000100000000000000000100001000000000000000001"; 
		when "0001" => Q <= "1000100000000000000000000010010000000000000000";
     	when "0010" => Q <= "0001010000000010000000000011000001000100000000";
		when "0011" => Q <= "0001110010101011000000000100001100010110000000";
		when "0100" => Q <= "0010010001000000000000010101000010000010000000";
		when "0101" => Q <= "0011000101010100100000001000111010101001000000";
		when "0110" => Q <= "0011010000010100110000000111000000000001010000";
		when "0111" => Q <= "0011110000000000100100001000000000000000000100";
		when "1000" => Q <= "0000100000000000000001001001000000101101100000";
		when "1001" => Q <= "0100110000100010101000001010000101010111001000";
		when "1010" => Q <= "0101010110001011000010000100100010000000000010";
		when others => Q <= "0000100000000000000000100001000000000000000001";
    	end case;	
end process;

end behavioral;
